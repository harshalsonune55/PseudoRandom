module xor2(
    input a,
    input b,
    output y
);
    assign y = a ^ b;
endmodule
